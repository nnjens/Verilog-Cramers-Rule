library verilog;
use verilog.vl_types.all;
entity cramer2 is
    port(
        HEX0            : out    vl_logic;
        HEX1            : out    vl_logic;
        HEX2            : out    vl_logic;
        HEX4            : out    vl_logic;
        HEX5            : out    vl_logic;
        HEX6            : out    vl_logic
    );
end cramer2;
